module mux_81_tb();
reg [8:0]i;
reg s0,s1,s2;
wire y;
mux_81 uut(.i(i),.s0(s0),.s1(s1),.s2(s2),.y(y));
initial 
begin
#100;s0=0;s1=0;s2=0;i[0]=1;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0;
#100;s0=0;s1=0;s2=1;i[0]=0;i[1]=1;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0;
#100;s0=0;s1=1;s2=0;i[0]=0;i[1]=0;i[2]=1;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=0;
#100;s0=0;s1=1;s2=1;i[0]=0;i[1]=0;i[2]=0;i[3]=1;i[4]=0;i[5]=0;i[6]=0;i[7]=0;
#100;s0=1;s1=0;s2=0;i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=1;i[5]=0;i[6]=0;i[7]=0;
#100;s0=1;s1=0;s2=1;i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=1;i[6]=0;i[7]=0;
#100;s0=1;s1=1;s2=0;i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=1;i[7]=0;
#100;s0=1;s1=1;s2=1;i[0]=0;i[1]=0;i[2]=0;i[3]=0;i[4]=0;i[5]=0;i[6]=0;i[7]=1;
end
endmodule
